// Dummy file to get SVUnit to run
